// `include "defines.v"

// module axi_rw # (
//     parameter RW_DATA_WIDTH     = 64,
//     parameter RW_ADDR_WIDTH     = 32,
//     parameter AXI_DATA_WIDTH    = 64,
//     parameter AXI_ADDR_WIDTH    = 32,
//     parameter AXI_ID_WIDTH      = 4,
//     parameter AXI_STRB_WIDTH    = AXI_DATA_WIDTH/8,
//     parameter AXI_USER_WIDTH    = 1
// )(
//     input                               clock,
//     input                               reset,

// 	input                               rw_valid_i,         //IF&MEM输入信号
// 	output                              rw_ready_o,         //IF&MEM输入信号
//     output reg [RW_DATA_WIDTH-1:0]      data_read_o,        //IF&MEM输入信号
//     input  [RW_DATA_WIDTH-1:0]          rw_w_data_i,        //IF&MEM输入信号
//     input  [RW_ADDR_WIDTH-1:0]          rw_addr_i,          //IF&MEM输入信号
//     input  [7:0]                        rw_size_i,          //IF&MEM输入信号



//     // Advanced eXtensible Interface
//     input                               axi_aw_ready_i,     //lite         
//     output                              axi_aw_valid_o,     //lite
//     output [AXI_ADDR_WIDTH-1:0]         axi_aw_addr_o,      //lite
//     output [2:0]                        axi_aw_prot_o,
//     output [AXI_ID_WIDTH-1:0]           axi_aw_id_o,
//     output [AXI_USER_WIDTH-1:0]         axi_aw_user_o,
//     output [7:0]                        axi_aw_len_o,       
//     output [2:0]                        axi_aw_size_o,
//     output [1:0]                        axi_aw_burst_o,
//     output                              axi_aw_lock_o,
//     output [3:0]                        axi_aw_cache_o,
//     output [3:0]                        axi_aw_qos_o,
//     output [3:0]                        axi_aw_region_o,

//     input                               axi_w_ready_i,      //lite              
//     output                              axi_w_valid_o,      //lite
//     output [AXI_DATA_WIDTH-1:0]         axi_w_data_o,       //lite
//     output [AXI_DATA_WIDTH/8-1:0]       axi_w_strb_o,       //lite
//     output                              axi_w_last_o,
//     output [AXI_USER_WIDTH-1:0]         axi_w_user_o,
    
//     output                              axi_b_ready_o,      //lite           
//     input                               axi_b_valid_i,      //lite
//     input  [1:0]                        axi_b_resp_i,       //lite            
//     input  [AXI_ID_WIDTH-1:0]           axi_b_id_i,
//     input  [AXI_USER_WIDTH-1:0]         axi_b_user_i,

//     input                               axi_ar_ready_i,     //lite              
//     output                              axi_ar_valid_o,     //lite
//     output [AXI_ADDR_WIDTH-1:0]         axi_ar_addr_o,      //lite
//     output [2:0]                        axi_ar_prot_o,
//     output [AXI_ID_WIDTH-1:0]           axi_ar_id_o,
//     output [AXI_USER_WIDTH-1:0]         axi_ar_user_o,
//     output [7:0]                        axi_ar_len_o,       //lite
//     output [2:0]                        axi_ar_size_o,      //lite
//     output [1:0]                        axi_ar_burst_o,
//     output                              axi_ar_lock_o,
//     output [3:0]                        axi_ar_cache_o,
//     output [3:0]                        axi_ar_qos_o,
//     output [3:0]                        axi_ar_region_o,
    
//     output                              axi_r_ready_o,      //lite            
//     input                               axi_r_valid_i,      //lite            
//     input  [1:0]                        axi_r_resp_i,
//     input  [AXI_DATA_WIDTH-1:0]         axi_r_data_i,       //lite
//     input                               axi_r_last_i,
//     input  [AXI_ID_WIDTH-1:0]           axi_r_id_i,
//     input  [AXI_USER_WIDTH-1:0]         axi_r_user_i
// );
    
//     // ------------------State Machine------------------TODO
    
//     // 写通道状态切换
    

//     // 读通道状态切换
    

//     // ------------------Write Transaction------------------
//     parameter AXI_SIZE      = $clog2(AXI_DATA_WIDTH / 8);
//     wire [AXI_ID_WIDTH-1:0] axi_id              = {AXI_ID_WIDTH{1'b0}};
//     wire [AXI_USER_WIDTH-1:0] axi_user          = {AXI_USER_WIDTH{1'b0}};
//     wire [7:0] axi_len      =  8'b0 ;
//     wire [2:0] axi_size     = AXI_SIZE[2:0];
//     // 写地址通道  以下没有备注初始化信号的都可能是你需要产生和用到的
//     assign axi_aw_valid_o   = w_state_addr;
//     assign axi_aw_addr_o    = rw_addr_i;
//     assign axi_aw_prot_o    = `AXI_PROT_UNPRIVILEGED_ACCESS | `AXI_PROT_SECURE_ACCESS | `AXI_PROT_DATA_ACCESS;  //初始化信号即可
//     assign axi_aw_id_o      = axi_id;                                                                           //初始化信号即可
//     assign axi_aw_user_o    = axi_user;                                                                         //初始化信号即可
//     assign axi_aw_len_o     = axi_len;
//     assign axi_aw_size_o    = axi_size;
//     assign axi_aw_burst_o   = `AXI_BURST_TYPE_INCR;                                                             
//     assign axi_aw_lock_o    = 1'b0;                                                                             //初始化信号即可
//     assign axi_aw_cache_o   = `AXI_AWCACHE_WRITE_BACK_READ_AND_WRITE_ALLOCATE;                                  //初始化信号即可
//     assign axi_aw_qos_o     = 4'h0;                                                                             //初始化信号即可
//     assign axi_aw_region_o  = 4'h0;                                                                             //初始化信号即可

//     // 写数据通道
//     assign axi_w_valid_o    = w_state_write;
//     assign axi_w_data_o     = rw_w_data_i ;
//     assign axi_w_strb_o     = rw_size_i;
//     assign axi_w_last_o     = 1'b0;
//     assign axi_w_user_o     = axi_user;                                                                         //初始化信号即可

//     // 写应答通道
//     assign axi_b_ready_o    = w_state_resp;

//     // ------------------Read Transaction------------------

//     // Read address channel signals
//     assign axi_ar_valid_o   = r_state_addr;
//     assign axi_ar_addr_o    = rw_addr_i;
//     assign axi_ar_prot_o    = `AXI_PROT_UNPRIVILEGED_ACCESS | `AXI_PROT_SECURE_ACCESS | `AXI_PROT_DATA_ACCESS;  //初始化信号即可
//     assign axi_ar_id_o      = axi_id;                                                                           //初始化信号即可                        
//     assign axi_ar_user_o    = axi_user;                                                                         //初始化信号即可
//     assign axi_ar_len_o     = axi_len;                                                                          
//     assign axi_ar_size_o    = axi_size;
//     assign axi_ar_burst_o   = `AXI_BURST_TYPE_INCR;
//     assign axi_ar_lock_o    = 1'b0;                                                                             //初始化信号即可
//     assign axi_ar_cache_o   = `AXI_ARCACHE_NORMAL_NON_CACHEABLE_NON_BUFFERABLE;                                 //初始化信号即可
//     assign axi_ar_qos_o     = 4'h0;                                                                             //初始化信号即可

//     // Read data channel signals
//     assign axi_r_ready_o    = r_state_read;

// endmodule