`include "defines.v"
module csr_reg (
    //TODO
);

endmodule //csr_reg