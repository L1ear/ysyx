// module icache(
//     input       
// );








// endmodule