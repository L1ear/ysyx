`include "defines.v"

module I_F (
);
    
endmodule