`include "defines.v"

module forwarding (
    
);

endmodule //forwarding