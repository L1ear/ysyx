module I_F (
);
    
endmodule