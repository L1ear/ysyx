module I_D (
    input                   instrc_i,

    output  [XLEN-1: 0]     rd;
    output  [XLEN-1: 0]     
);
    
endmodule